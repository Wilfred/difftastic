architecture a of e is
begin
end architecture b;
              -- ^ error.misspeling.name
