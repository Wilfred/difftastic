package pkg is
end package foo;
         -- ^ error.misspeling.name

