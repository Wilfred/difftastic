entity ent is
end entity foo;
        -- ^ error.misspeling.name
