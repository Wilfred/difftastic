package body pkg is
end package body foo;
              -- ^ error.misspeling.name

